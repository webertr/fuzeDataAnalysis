*
* This circuit contains a capacitor and an inductor with
* is designed to simulate the fuze circuit
*

* Global parameters for simulation
*.param corn=2


************************************************************************************************
* Thyristor Bank
************************************************************************************************

* Instance of capacitor and thyristor switch
xthyBank1 1 0 r1p r1n id1 it1p it1n vthyBank 
          +trigTime1a=10u trigTime1b=11u
          +initialVoltage=7k
	  +capValue=830u

* Instance of capacitor and thyristor switch
xthyBank2 1 0 r2p r2n id2 it2p it2n vthyBank 
          +trigTime1a=10u trigTime1b=11u
          +initialVoltage=7k
	  +capValue=830u

* Instance of capacitor and thyristor switch
xthyBank3 1 0 r3p r3n id3 it3p it3n vthyBank 
          +trigTime1a=10u trigTime1b=11u
          +initialVoltage=7k
	  +capValue=830u

* Instance of capacitor and thyristor switch
xthyBank4 1 0 r4p r4n id4 it4p it4n vthyBank 
          +trigTime1a=10u trigTime1b=11u
          +initialVoltage=7k
	  +capValue=830u

* Instance of capacitor and thyristor switch
xthyBank5 1 0 r5p r5n id5 it5p it5n vthyBank 
          +trigTime1a=10u trigTime1b=11u
          +initialVoltage=7k
	  +capValue=830u

* Instance of capacitor and thyristor switch
xthyBank6 1 0 r6p r6n id6 it6p it6n vthyBank 
          +trigTime1a=10u trigTime1b=11u
          +initialVoltage=7k
	  +capValue=830u

* Instance of capacitor and thyristor switch
xthyBank7 1 0 r7p r7n id7 it7p it7n vthyBank 
          +trigTime1a=10u trigTime1b=11u
          +initialVoltage=7k
	  +capValue=830u

* Instance of capacitor and thyristor switch
xthyBank8 1 0 r8p r8n id8 it8p it8n vthyBank 
          +trigTime1a=10u trigTime1b=11u
          +initialVoltage=7k
	  +capValue=830u

* Instance of capacitor and thyristor switch
xthyBank9 1 0 r9p r9n id9 it9p it9n vthyBank 
          +trigTime1a=10u trigTime1b=11u
          +initialVoltage=7k
	  +capValue=830u

* Instance of capacitor and thyristor switch
xthyBank10 1 0 r10p r10n id10 it10p it10n vthyBank 
          +trigTime1a=10u trigTime1b=11u
          +initialVoltage=7k
	  +capValue=830u

* Instance of capacitor and thyristor switch
xthyBank11 1 0 r11p r11n id11 it11p it11n vthyBank 
          +trigTime1a=10u trigTime1b=11u
          +initialVoltage=7k
	  +capValue=830u

* Instance of capacitor and thyristor switch
xthyBank12 1 0 r12p r12n id12 it12p it12n vthyBank 
          +trigTime1a=10u trigTime1b=11u
          +initialVoltage=7k
	  +capValue=830u


************************************************************************************************
* Ignitron Bank
************************************************************************************************

* Instance of ignitron bank module
xignBank1 1 0 ri1p ri1n rtot1p rtot1n rs1p rs1n capv1 vignBank 
          +trigTime1a=10u trigTime1b=11u
          +initialVoltage=7k
	  +capValue=37u

* Instance of ignitron bank module
xignBank2 1 0 ri2p ri2n rtot2p rtot2n rs2p rs2n capv2 vignBank 
          +trigTime1a=10u trigTime1b=11u
          +initialVoltage=7k
	  +capValue=37u

* Instance of ignitron bank module
xignBank3 1 0 ri3p ri3n rtot3p rtot1n rs3p rs3n capv3 vignBank 
          +trigTime1a=10u trigTime1b=11u
          +initialVoltage=7k
	  +capValue=37u

* Instance of ignitron bank module
xignBank4 1 0 ri4p ri4n rtot4p rtot4n rs4p rs4n capv4 vignBank 
          +trigTime1a=10u trigTime1b=11u
          +initialVoltage=7k
	  +capValue=37u

* Instance of ignitron bank module
xignBank5 1 0 ri5p ri5n rtot5p rtot5n rs5p rs5n capv5 vignBank 
          +trigTime1a=10u trigTime1b=11u
          +initialVoltage=7k
	  +capValue=37u

* Instance of ignitron bank module
xignBank6 1 0 ri6p ri6n rtot6p rtot6n rs6p rs6n capv6 vignBank 
          +trigTime1a=10u trigTime1b=11u
          +initialVoltage=7k
	  +capValue=37u


************************************************************************************************
* Bank load
************************************************************************************************

* Shunt resistance
RS 1 2 1u

* Plasma impedance
xplasmaLoad1 2 0 vplasmaload

* Snubber impedance
xsnubberLoad1 2 0 vsnubber

* Dummy load
xdummyLoad1 2 0 vdummyload



************************************************************************************************
* Ignitron bank module model
************************************************************************************************

* Model of a capacitor and ignitron bank module.
.subckt vignBank 11 10 2 3 7 8 12 13 1
                 +trigTime1a=0.3 trigTime1b=0.31
                 +initialVoltage=5k
		 +capValue=37u

* 10 = the ground. Ignitron = NL8900
C1 1 10 capValue ic=initialVoltage
L1 1 2 10n
R1 2 3 6.3m
L2 3 4 120n
R2 4 5 0.1m
SwitchOUT 5 6 99 10 switch_out off 
L3 6 7 500n
R3 7 8 1.9m
L4 8 11 640n
SwitchCB 3 9 3 10 switch_cb on
L5 9 12 130n
RS 12 13 1u
R4 13 10 0.1m

* Ignitron switch model control voltage
v1 99 10 DC PWL(0 0 trigTime1a 0 trigTime1b 1)

* Models
* Switch model for output
* vt = on threshold, vh = hystersis, ron = on resistance
* roff = off resistance
.model switch_out sw vt=1.0 vh=0 ron=0.1m roff=1gig

* Switch model for cb
* vt = on threshold, vh = hystersis, ron = on resistance
* roff = off resistance The switch trips at (Vt − Vh) and (Vt + Vh)
.model switch_cb sw vt=5000 vh=5000 ron=1gig roff=0.1m

.ends




************************************************************************************************
* Thyristor bank module model
************************************************************************************************

* Model of a capacitor and thyristor switch.
.subckt vthyBank 14 10 1 2 33 11 12
                 +trigTime1a=0.3 trigTime1b=0.31
                 +initialVoltage=5k
		 +capValue=840u

* 10 = the ground
C1 1 10 capValue ic=initialVoltage
R41 1 2 1m
L35 2 3 40n
L3 3 4 200n
R7 4 5 6m
diode0 33 5 DCLAMP
RS 33 10 1u
C11 5 6 1u ic=initialVoltage
R10 6 10 4
switch1 5 8 99 10 switch1 off 
diode6 8 9 DCLAMP
L23 9 11 200n
R11 11 12 3.33m
L10 12 13 1.122u
L47 13 14 300n

* Thyristor switch model control voltage
v1 99 10 DC PWL(0 0 trigTime1a 0 trigTime1b 1)
* Models
* Switch model
* vt = on threshold, vh = hystersis, ron = on resistance
* roff = off resistance
.model switch1 sw vt=0.1 vh=0 ron=0.5m roff=1gig
* Diode model
* DC Parameters:
* BV = Reverse breakdown voltage, IBV = Current at breakdown voltage
* IK = Forward Knee Current, IKR = Reverse Knee Current
* IS = Saturation Current (Scaled by "AREA" in instance declaration)
* JSW = Side wall saturation, N = Emission Coefficient
* RS = Ohmic resistance
.model DCLAMP D rs=0.17m

.ends



************************************************************************************************
* Module of snubbers
************************************************************************************************

* Model of the snubbers used on the FuZE experiment
.subckt vsnubber 1 4
                 +resValue=0.07
		 +capValue=0.6u
		 +inductValue=25n

* Snubber inductance
L1 1 2 inductValue
* Snubber capacitor
C1 2 3 capValue
* Snubber resistance
R1 3 4 resValue

.ends



************************************************************************************************
* Model of dummy load
************************************************************************************************

* Model of the dummy load used on the FuZE experiment
.subckt vdummyload 1 3
                 +resValue=1.7
		 +inductValue=5u

* Dummy inductance
L1 1 2 inductValue
* Dummy resistance
R1 2 3 resValue

.ends


************************************************************************************************
* Model of plasma load
************************************************************************************************

* Model of the plasma load used on the FuZE experiment
.subckt vplasmaload 1 3
                 +resValue=5m
		 +inductValue=152n

* Plasma resistance
R1 1 2 resValue
* Plasma inductance
L1 2 3 inductValue

.ends



* Starting control statements
.control

* Setting output file type
set filetype=ascii
* Specifying time domain to solve solution for and enabling I.C.'s
*.tran tstep tstop <tstart <tmax>> <uic>
* tstep = suggested step time, tstop = stop time
* tstart = start time (defaults to 0)
* tmax = maximum time step, uic = use initial conditions
tran 5n 500u 0 50n uic
* Plotting 
*plot v(5)
* Writting output file for I from Ignitron bank Capacitor
write ic1.txt (v(ri1p)-v(ri1n))/6.3m/1000
* Writting output file for total ip
write ip.txt (v(1)-v(2))/1u/1000
* Writting output file for ignitron out 1
write iout1.txt (v(rtot1p)-v(rtot1n))/1.9m/1000
* Writting output file for ignitron cb 1
write icb1.txt (v(rs1n)-v(rs1p))/1u/1000
* Writting output for vgap
write vgap.txt v(2)/1000
* Writting voltage at ignitron cb
write vigcb.txt v(ri1n)/1000
* Writting voltage from ignitron capacitor 1
write vcap1.txt v(capv1)/1000
* Writting voltage from ignitron capacitor 1
write vtcap1.txt v(r1p)/1000

* Ending control statement
.endc

* Ending circuit simulation
.end