*
* This circuit contains a capacitor and an inductor with
* is designed to simulate the fuze circuit
*

* Global parameters for simulation
*.param corn=2

* Instance of ignitron bank module
xignBank1 1 0 r1p r1n r4p r3p r3n vignBank 
          +trigTime1a=10u trigTime1b=11u
          +initialVoltage=5k
	  +capValue=37u

* Shunt resistance
RS 1 2 1u

* Plasma impedance
xplasmaLoad1 2 0 vplasmaload

* Snubber impedance
xsnubberLoad1 2 0 vsnubber

* Dummy load
xdummyLoad1 2 0 vdummyload



* Model of a capacitor and ignitron bank module.
.subckt vignBank 11 10 2 3 12 7 8
                 +trigTime1a=0.3 trigTime1b=0.31
                 +initialVoltage=5k
		 +capValue=37u

* 10 = the ground. Ignitron = NL8900
C1 1 10 capValue ic=initialVoltage
L1 1 2 10n
R1 2 3 6.3m
L2 3 4 120n
R2 4 5 0.1m
SwitchOUT 5 6 99 10 switch_out off 
L3 6 7 500n
R3 7 8 1.9m
L4 8 11 640n
SwitchCB 3 9 3 10 switch_cb on
L5 9 12 130n
R4 12 10 0.1m

* Ignitron switch model control voltage
v1 99 10 DC PWL(0 0 trigTime1a 0 trigTime1b 1)

* Models
* Switch model for output
* vt = on threshold, vh = hystersis, ron = on resistance
* roff = off resistance
.model switch_out sw vt=1.0 vh=0 ron=0.1m roff=1gig

* Switch model for cb
* vt = on threshold, vh = hystersis, ron = on resistance
* roff = off resistance
.model switch_cb sw vt=5000 vh=5000 ron=1gig roff=0.1m

.ends

* Model of the snubbers used on the FuZE experiment
.subckt vsnubber 1 4
                 +resValue=0.07
		 +capValue=0.6u
		 +inductValue=25n

* Snubber inductance
L1 1 2 inductValue
* Snubber capacitor
C1 2 3 capValue
* Snubber resistance
R1 3 4 resValue

.ends

* Model of the dummy load used on the FuZE experiment
.subckt vdummyload 1 3
                 +resValue=1.7
		 +inductValue=5u

* Dummy inductance
L1 1 2 inductValue
* Dummy resistance
R1 2 3 resValue

.ends

* Model of the plasma load used on the FuZE experiment
.subckt vplasmaload 1 3
                 +resValue=5m
		 +inductValue=152n

* Plasma resistance
R1 1 2 resValue
* Plasma inductance
L1 2 3 inductValue

.ends


* Starting control statements
.control

* Setting output file type
set filetype=ascii
* Specifying time domain to solve solution for and enabling I.C.'s
*.tran tstep tstop <tstart <tmax>> <uic>
* tstep = suggested step time, tstop = stop time
* tstart = start time (defaults to 0)
* tmax = maximum time step, uic = use initial conditions
tran 5n 500u 0 50n uic
* Plotting 
*plot v(5)
* Writting output file for I from Capacitor
write ic1.txt (v(r1p)-v(r1n))/6.3m/1000
* Writting output file for total ip
write ip.txt (v(1)-v(2))/1u/1000
* Writting output file for ignitron out 1
write iout1.txt (v(r3p)-v(r3n))/1.9m/1000
* Writting output file for ignitron cb 1
write icb1.txt (v(r4p)-v(0))/0.1m/1000
* Writting output for vgap
write vgap.txt v(2)/1000

* Ending control statement
.endc

* Ending circuit simulation
.end